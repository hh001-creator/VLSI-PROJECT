.include "TSMC_180nm.txt"
.include "logicgates.cir"
.param LAMBDA = 0.09u
.param width_N = {10*LAMBDA}
.param width_P = {2*width_N}
.param SUPPLY = 1.8
.global gnd vdd

VDD vdd gnd 1.8
**INPUTS**
Vin1 A1 gnd pulse(0 1.8 0 0 0 100ns 0)
Vin2 A2 gnd pulse(0 1.8 0 0 0 100ns 0)
Vin3 A3 gnd pulse(0 1.8 0 0 0 100ns 0)
Vin4 A4 gnd pulse(0 1.8 0 0 0 100ns 0)

Vin5 B1 gnd pulse(0 1.8 0 0 0 100ns 0)
Vin6 B2 gnd pulse(0 1.8 0 0 0 100ns 0)
Vin7 B3 gnd pulse(0 1.8 0 0 0 100ns 0)
Vin8 B4 gnd pulse(0 1.8 0 0 0 100ns 0) 



.subckt cla ina1 ina2 ina3 ina4 inb1 inb2 inb3 inb4 out1 out2 out3 out4 out5 hi lo
*P1 P2 P3 P4
xX1 P1 ina1 inb1 hi lo cmosxor
xX2 P2 ina2 inb2 hi lo cmosxor
xX3 P3 ina3 inb3 hi lo cmosxor
xX4 P4 ina4 inb4 hi lo cmosxor

** G1 G2 G3 G4
xA1 G1 ina1 inb1 hi lo cmosand
xA2 G2 ina2 inb2 hi lo cmosand
xA3 G3 ina3 inb3 hi lo cmosand
xA4 G4 ina4 inb4 hi lo cmosand

** C1 = 0 
** C2 = G1
** C3 = G2 + P2G1
**Op1 = P2G1
xAn1 Op1 P2 G1 hi lo cmosand
xO1 C3 G2 Op1 hi lo cmosor

**C4 = G3 + P3G2 + P3P2G1
** Op2 = P3G2
xAn2 Op2 P3 G2 hi lo cmosand
** Op3 = P3P2G1
xAn3 Op3 P3 Op1 hi lo cmosand
**Op4 =  G3 + P3G2
xO2 Op4 G3 Op2 hi lo cmosor
** C4 = Op4 + Op3
xO3 C4 Op4 Op3 hi lo cmosor

** C5 = G4 + P4G3 + P4P3G2 + P4P3P2G1 = G4 + ot1 + ot2  + ot3
** Ot1 = P4G3
xAnd1 Ot1 P4 G3 hi lo cmosand
** Ot2 = P4P3G2
xAnd2 Ot2 P4 Op2 hi lo cmosand
** Ot3 = P4P3P2G1
xAnd3 Ot3 P4 Op4 hi lo cmosand
** Ot4 = G4 + Ot1
xOrg1 Ot4 G4 Ot1 hi lo cmosor
** Ot5 = Ot2 + Ot3
xOrg2 Ot5 Ot2 Ot3 hi lo cmosor
** out5 = Ot4 + Ot5 => Cout
xOrg3 out5 Ot5 Ot4 hi lo cmosor

xXo1 out1 P1 lo hi lo cmosxor
xXo2 out2 P2 G1 hi lo cmosxor
xXo3 out3 P3 C3 hi lo cmosxor
xXo4 out4 P4 C4 hi lo cmosxor

.ends cla


xcla1 A1 A2 A3 A4 B1 B2 B3 B4 S1 S2 S3 S4 Cout vdd gnd cla 
.tran 10ps 50ns 

*.measure tran tplh
*+ TRIG v(A) VAL = 'SUPPLY/2' FALL = 1
*+ TARG V(OpAnd) VAL = 'SUPPLY/2' RISE = 1
*.measure tran tphl
*+ TRIG V(A) VAL = 'SUPPLY/2' RISE = 1
*+ TARG V(OpAnd) VAL = 'SUPPLY/2' FALL = 1

.control
	run
	set hcopypscolor = 1
	set color0 = white
	set color1 = black
	
.endc
.end
