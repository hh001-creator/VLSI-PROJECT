
.include "TSMC_180nm.txt"
.include "cmoslogic.cir"
.include "logicgates.cir"
.include "cla.cir"
.include "Dff.cir"

.param LAMBDA = 0.09u
.param width_N = {10*LAMBDA}
.param width_P = {2*width_N}
.param SUPPLY = 1.8
.global gnd vdd

VDD vdd gnd 1.8
**INPUTS**
Vin1 A1 gnd pulse(0 1.8 0 0 0 100ns 0)
Vin2 A2 gnd pulse(0 1.8 0 0 0 100ns 0)
Vin3 A3 gnd pulse(0 1.8 0 0 0 100ns 0)
Vin4 A4 gnd pulse(0 1.8 0 0 0 100ns 0)

Vin5 B1 gnd pulse(0 1.8 0 0 0 100ns 0)
Vin6 B2 gnd pulse(0 1.8 0 0 0 100ns 0)
Vin7 B3 gnd pulse(0 1.8 0 0 0 100ns 0)
Vin8 B4 gnd pulse(0 1.8 0 0 0 100ns 0) 

Vin9 clk     gnd pulse( 0 1.8 0.2ns 0ps 0ps 0.2ns 0.4ns 0 )
Vin10 clk_bar gnd pulse( 1.8 0 0.2ns 0ps 0ps 0.2ns 0.4ns 0 )

xDff1 O1 A1 clk clk_bar vdd gnd DFlipFlop 
xDff2 O2 A2 clk clk_bar vdd gnd DFlipFlop
xDff3 O3 A3 clk clk_bar vdd gnd DFlipFlop
xDff4 O4 A4 clk clk_bar vdd gnd DFlipFlop

xDff5 O5 B1 clk clk_bar vdd gnd DFlipFlop
xDff6 O6 B2 clk clk_bar vdd gnd DFlipFlop
xDff7 O7 B3 clk clk_bar vdd gnd DFlipFlop
xDff8 O8 B4 clk clk_bar vdd gnd DFlipFlop

xCLA O1 O2 O3 O4 O5 O6 O7 O8 SP1 SP2 SP3 SP4 CO vdd gnd cla

xDf1 S1 SP1 clk clk_bar vdd gnd DFlipFlop
xDf2 S2 SP2 clk clk_bar vdd gnd DFlipFlop
xDf3 S3 SP3 clk clk_bar vdd gnd DFlipFlop
xDf4 S4 SP4 clk clk_bar vdd gnd DFlipFlop

xDf5 Cout CO clk clk_bar vdd gnd DFlipFlop  


.tran 20ps 100ns 


.control
	run
	set hcopypscolor = 1
	set color0 = white
	set color1 = black
	
.endc
.end
