And Gate Using Transmission Gate
.include "TSMC_180nm.txt"
.param LAMBDA = 0.09u
.param width_N = {10*LAMBDA}
.param width_P = {2*width_N}
.param SUPPLY = 1.8
.global gnd vdd

Vin1 A gnd pulse(0 1.8 20ns 0 0 50ns 0)
Vin2 B gnd pulse(0 1.8 30ns 0 0 50ns 0)

.subckt cmosinv out in hi lo 
M1 out in lo lo 
+ CMOSN W={width_N} L={2*LAMBDA} 
+ AS={5*width_N*LAMBDA} PS={10*LAMBDA+2*width_N} 
+ AD={5*width_N*LAMBDA} PD={10*LAMBDA+2*width_N}

M2 out in hi hi 
+ CMOSP W={width_P} L={2*LAMBDA} 
+ AS={5*width_P*LAMBDA} PS={10*LAMBDA+2*width_P} 
+ AD={5*width_P*LAMBDA} PD={10*LAMBDA+2*width_P}

.ends cmosinv

.subckt TG out in1 in2 in3 hi lo
M1 out in3 in1 hi
+ CMOSP W={width_P} L={2*LAMBDA} 
+ AS={5*width_P*LAMBDA} PS={10*LAMBDA+2*width_P} 
+ AD={5*width_P*LAMBDA} PD={10*LAMBDA+2*width_P}

M2 out in2 in1 hi
+ CMOSN W={width_N} L={2*LAMBDA} 
+ AS={5*width_N*LAMBDA} PS={10*LAMBDA+2*width_N} 
+ AD={5*width_N*LAMBDA} PD={10*LAMBDA+2*width_N}

.ends TG

.subckt cmosxor out in1 in2 hi lo
xI1 in1_bar in1 hi lo cmosinv
xI2 in2_bar in2 hi lo cmosinv

xTG1 out in1 in2_bar in2 hi lo TG
xTG2 out in1_bar in2 in2_bar hi lo TG 
.ends cmosxor

xA1 out A B vdd gnd cmosxor
.tran 10ps 50ns 

.control
	run
    set hcopypscolor = 1
	set color0 = white
	set color1 = black
.endc

.end