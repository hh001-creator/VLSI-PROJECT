.include TSMC_180nm.txt
.param LAMBDA = 0.09u
.param width_N = {10*LAMBDA}
.param width_P = {2*width_N}
.param SUPPLY = 1.8
.global gnd vdd

VDD vdd gnd 1.8
**INPUTS**
Vin1 A1 gnd pulse(0 1.8 0 0 0 100ns 0)
Vin2 A2 gnd pulse(0 1.8 0 0 0 100ns 0)
Vin3 A3 gnd pulse(0 1.8 0 0 0 100ns 0)
Vin4 A4 gnd pulse(0 1.8 0 0 0 100ns 0)

Vin5 B1 gnd pulse(0 1.8 5ns 0 0 100ns 0)
Vin6 B2 gnd pulse(0 0 0 0 0 100ns 0)
Vin7 B3 gnd pulse(0 0 0 0 0 100ns 0)
Vin8 B4 gnd pulse(0 0 0 0 0 100ns 0) 

.subckt cmosinv out in hi lo 
M1 out in lo lo 
+ CMOSN W={width_N} L={2*LAMBDA} 
+ AS={5*width_N*LAMBDA} PS={10*LAMBDA+2*width_N} 
+ AD={5*width_N*LAMBDA} PD={10*LAMBDA+2*width_N}

M2 out in hi hi 
+ CMOSP W={width_P} L={2*LAMBDA} 
+ AS={5*width_P*LAMBDA} PS={10*LAMBDA+2*width_P} 
+ AD={5*width_P*LAMBDA} PD={10*LAMBDA+2*width_P}

.ends cmosinv

.subckt cmosnand out in1 in2 hi lo
M1 out in1 hi hi 
+ CMOSP W={width_P} L={2*LAMBDA} 
+ AS={5*width_P*LAMBDA} PS={10*LAMBDA+2*width_P} 
+ AD={5*width_P*LAMBDA} PD={10*LAMBDA+2*width_P}

M2 out in2 hi hi
+ CMOSP W={width_P} L={2*LAMBDA} 
+ AS={5*width_P*LAMBDA} PS={10*LAMBDA+2*width_P} 
+ AD={5*width_P*LAMBDA} PD={10*LAMBDA+2*width_P}

M3 out in1 C gnd
+ CMOSN W={width_N} L={2*LAMBDA} 
+ AS={5*width_N*LAMBDA} PS={10*LAMBDA+2*width_N} 
+ AD={5*width_N*LAMBDA} PD={10*LAMBDA+2*width_N}

M4 C in2 gnd gnd
+ CMOSN W={width_N} L={2*LAMBDA} 
+ AS={5*width_N*LAMBDA} PS={10*LAMBDA+2*width_N} 
+ AD={5*width_N*LAMBDA} PD={10*LAMBDA+2*width_N}

.ends cmosnand

************AND GATE************

.subckt cmosand out in1 in2 hi lo
xND1 out1 in1 in2 hi lo cmosnand
xI1 out out1 hi lo cmosinv
.ends cmosand
*******************************

************OR GATE************
.subckt cmosor out in1 in2 hi lo
xI2 o1 in1 hi lo cmosinv
xI3 o2 in2 hi lo cmosinv
xND2 out o1 o2 vdd gnd cmosnand
.ends cmosor

*******************************

************XOR GATE************
.subckt cmosxor out in1 in2 hi lo
xND3 o1 in1 in2 vdd gnd cmosnand
xND4 o2 in1 o1 vdd gnd cmosnand
xND5 o3 o1 in2 vdd gnd cmosnand
xND6 out o2 o3 vdd gnd cmosnand
.ends cmosxor
*******************************

xX1 P1 A1 B1 vdd gnd cmosxor
xX2 P2 A2 B2 vdd gnd cmosxor
xX3 P3 A3 B3 vdd gnd cmosxor
xX4 P4 A4 B4 vdd gnd cmosxor

xA1 G1 A1 B1 vdd gnd cmosand
xA2 G2 A2 B2 vdd gnd cmosand
xA3 G3 A3 B3 vdd gnd cmosand
xA4 G4 A4 B4 vdd gnd cmosand

**********C3******************
xAn1 Op1 P2 G1 vdd gnd cmosand
xO1 C3 G2 Op1 vdd gnd cmosor
******************************

xAn2 Op2 P3 G2 vdd gnd cmosand

**********P3P2G1***************
xAn3 Op3 P3 P2 vdd gnd cmosand
xAn4 Op4 Op3 G1 vdd gnd cmosand
********************************
*********G3 + P3G2*************
xO2 Op5 G3 Op2 vdd gnd cmosor
*******************************

**************C4***************
xO3 C4 Op5 Op4 vdd gnd cmosor
******************************

xAn5 Op6 P4 C4 vdd gnd cmosand
xO4 C5 G4 Op6 vdd gnd cmosor

xXo1 S1 P1 gnd vdd gnd cmosxor
xXo2 S2 P2 G1 vdd gnd cmosxor
xXo3 S3 P3 C3 vdd gnd cmosxor
xXo4 S4 P4 C4 vdd gnd cmosxor
.tran 10ps 50ns 

*.measure tran tplh
*+ TRIG v(A) VAL = 'SUPPLY/2' FALL = 1
*+ TARG V(OpAnd) VAL = 'SUPPLY/2' RISE = 1
*.measure tran tphl
*+ TRIG V(A) VAL = 'SUPPLY/2' RISE = 1
*+ TARG V(OpAnd) VAL = 'SUPPLY/2' FALL = 1

.control
	run
	set hcopypscolor = 1
	set color0 = white
	set color1 = black
	
.endc
.end
